library ieee;
    use ieee.std_logic_1164.all;

entity carry_save_tree_adder is
    generic (
        N_BITS          : POSITIVE; -- Number of bits per addend
        N_INPUTS        : POSITIVE; -- Number of addends
        TWOS_COMPLEMENT : BOOLEAN   -- Use 2's complement extension
    );

    port (
        addends : in    STD_LOGIC_VECTOR(N_BITS * N_INPUTS - 1 downto 0); -- Inputs: addends concatenated
        sum     : out   STD_LOGIC_VECTOR(N_BITS + N_INPUTS - 1 downto 0)  -- Outputs
    );
end entity carry_save_tree_adder;

architecture behavioral of carry_save_tree_adder is
    -- Constants
    constant TOT_CSA_N : POSITIVE := N_INPUTS - 2; -- Total number of carry save adders of the tree

    -- Level map
    type level_map_type is array (0 to TOT_CSA_N - 1) of INTEGER; -- Array of levels for each carry save adder
    -- Compute the levels of each carry save adder
    function compute_levels (
        n_in  : POSITIVE;                  -- Number of inputs
        n_csa : POSITIVE                   -- Number of carry save adders
    ) return level_map_type is
        variable map_arr : level_map_type; -- Return value

        variable w       : INTEGER;  -- Number of wires of the current level
        variable new_csa : INTEGER;  -- Number of carry save adders of the current level
        variable l       : POSITIVE; -- Current level
    begin
        w       := n_in;             -- First level has number of wires equal to number of inputs
        new_csa := 0;                -- No carry save adders at the beginning
        l       := 1;                -- Start at level 1
        -- Loop over each carry save adder
        for i in 0 to n_csa - 1 loop
            -- Check if the current level is full
            if (w <= 2) then
                w       := w + (new_csa * 2); -- Set the new number of wires for the next level
                new_csa := 0;                 -- Reset the number of carry save adders for the next level
                l       := l + 1;             -- Increment the level
            end if;

            map_arr(i) := l; -- Set the level of the current carry save adder

            w       := w - 3;       -- Consume 3 wires
            new_csa := new_csa + 1; -- Increment the number of carry save adders of the current level
        end loop;

        return map_arr;
    end function compute_levels;

    constant CSA_LEVELS : level_map_type := compute_levels(N_INPUTS, TOT_CSA_N); -- Levels of each carry save adder

    -- Signals for recursive assignment
    -- Compute the size of the added signals resulting from each carry save adder
    function compute_signal_sizes (
        n_bits    : POSITIVE;      -- Number of bits of the inputs
        level_map : level_map_type -- Levels of each carry save adder
    ) return INTEGER is
        variable size : INTEGER;   -- Return value
    begin
        size := 0;                 -- Initialize the return value to 0

        -- Loop over each carry save adder
        for i in 0 to level_map'length - 1 loop
            -- The size of each output of a carry save adder is equal to `n_bits + csa_level` (the level start from 1)
            -- Each carry save adder has 2 outputs
            size := size + (n_bits + level_map(i)) * 2;
        end loop;

        return size;
    end function compute_signal_sizes;

    constant SIGNAL_SIZES : INTEGER := compute_signal_sizes(N_BITS, CSA_LEVELS); -- Size of the added signals
    -- Total size of the structure that contains the inputs and the added signals generated by the carry save adders
    constant TOT_SIGNALS_N : POSITIVE := N_INPUTS * N_BITS + SIGNAL_SIZES;
    constant TOT_WIRES_N   : POSITIVE := N_INPUTS + 2 * TOT_CSA_N; -- Total number of wires

    -- Recursive assignment signals structure
    signal recursive_signals : STD_LOGIC_VECTOR(TOT_SIGNALS_N - 1 downto 0);

    -- Signal offsets
    type int_array is array (0 to TOT_WIRES_N - 1) of INTEGER;
    -- Compute the offset of each wire
    function compute_wire_offset (
        n_bits_in : POSITIVE;              -- Number of bits of the inputs
        n_in      : POSITIVE;              -- Number of inputs
        lvl_map   : level_map_type         -- Levels of each carry save adder
    ) return int_array is
        variable offsets      : int_array; -- Return value
        variable current_pos  : INTEGER;   -- Current offset position
        variable signal_width : INTEGER;   -- Width of the current signal
    begin
        current_pos := 0;                  -- Current offset position

        -- Offset of the inputs signals
        for i in 0 to n_in - 1 loop
            offsets(i)  := current_pos;
            current_pos := current_pos + n_bits_in; -- Update the current offset position with the width of the input
        end loop;

        -- Offset of the carry save adder result signals
        for k in 0 to lvl_map'length - 1 loop
            -- The width of the output signal of a carry save adder is equal to `n_bits_in + csa_level`
            -- (starting from level 1)
            signal_width := n_bits_in + lvl_map(k);

            -- PS output
            offsets(n_in + k * 2) := current_pos;
            current_pos           := current_pos + signal_width;

            -- CV output
            offsets(n_in + k * 2 + 1) := current_pos;
            current_pos               := current_pos + signal_width;
        end loop;

        return offsets;
    end function compute_wire_offset;

    -- List of the offsets of each wire
    constant WIRE_OFFSETS : int_array := compute_wire_offset(N_BITS, N_INPUTS, CSA_LEVELS);

    -- Components
    component carry_save_adder is
        generic (
            N : POSITIVE
        );

        port (
            a, b, c : in    STD_LOGIC_VECTOR(n - 1 downto 0);
            ps, cv  : out   STD_LOGIC_VECTOR(n - 1 downto 0)
        );
    end component carry_save_adder;

    component extender is
        generic (
            N_IN            : POSITIVE;
            N_OUT           : POSITIVE;
            TWOS_COMPLEMENT : BOOLEAN
        );

        port (
            data_in  : in    STD_LOGIC_VECTOR(N_IN - 1 downto 0);
            data_out : out   STD_LOGIC_VECTOR(N_OUT - 1 downto 0)
        );
    end component extender;

    component ripple_carry_adder is
        generic (
            N : POSITIVE
        );

        port (
            a, b : in    STD_LOGIC_VECTOR(n - 1 downto 0);
            cin  : in    STD_LOGIC;
            s    : out   STD_LOGIC_VECTOR(n - 1 downto 0);
            cout : out   STD_LOGIC
        );
    end component ripple_carry_adder;

begin
    -- Setting the inputs in the recursive assignment structure
    recursive_signals(N_BITS * N_INPUTS - 1 downto 0) <= addends;

    -- Instantiating of each carry save adder
    csa: for i in 0 to TOT_CSA_N - 1 generate
        -- Level
        constant LVL : INTEGER := CSA_LEVELS(i); -- Level of the current carry save adder (starting from 1)
        -- Current signal width
        constant CURRENT_CSA_WIDTH : POSITIVE := N_BITS + LVL - 1; -- Width of the current carry save adder

        -- Indexes
        -- Inputs
        constant IDX_A : INTEGER := i * 3;
        constant IDX_B : INTEGER := i * 3 + 1;
        constant IDX_C : INTEGER := i * 3 + 2;
        -- Outputs
        constant IDX_PS : INTEGER := N_INPUTS + i * 2;
        constant IDX_CV : INTEGER := N_INPUTS + i * 2 + 1;

        -- Signals
        signal a_i, b_i, c_i : STD_LOGIC_VECTOR(CURRENT_CSA_WIDTH - 1 downto 0);
        signal ps_i, cv_i    : STD_LOGIC_VECTOR(CURRENT_CSA_WIDTH - 1 downto 0);
    begin
        -- Extending the inputs
        -- Extending applied only if the signal comes form a earlier layer that the previous one
        -- If the signal comes from a later layer, it will apply an extension of 0 (ignored by the compiler)
        ext_a: component extender
            generic map (
                N_IN            => (WIRE_OFFSETS(IDX_A + 1) - WIRE_OFFSETS(IDX_A)),
                N_OUT           => CURRENT_CSA_WIDTH,
                TWOS_COMPLEMENT => TWOS_COMPLEMENT
            )

            port map (
                data_in  => recursive_signals(WIRE_OFFSETS(IDX_A + 1) - 1 downto WIRE_OFFSETS(IDX_A)),
                data_out => a_i
            );
        ext_b: component extender
            generic map (
                N_IN            => (WIRE_OFFSETS(IDX_B + 1) - WIRE_OFFSETS(IDX_B)),
                N_OUT           => CURRENT_CSA_WIDTH,
                TWOS_COMPLEMENT => TWOS_COMPLEMENT
            )

            port map (
                data_in  => recursive_signals(WIRE_OFFSETS(IDX_B + 1) - 1 downto WIRE_OFFSETS(IDX_B)),
                data_out => b_i
            );
        ext_c: component extender
            generic map (
                N_IN            => (WIRE_OFFSETS(IDX_C + 1) - WIRE_OFFSETS(IDX_C)),
                N_OUT           => CURRENT_CSA_WIDTH,
                TWOS_COMPLEMENT => TWOS_COMPLEMENT
            )

            port map (
                data_in  => recursive_signals(WIRE_OFFSETS(IDX_C + 1) - 1 downto WIRE_OFFSETS(IDX_C)),
                data_out => c_i
            );

        -- Instantiating of the carry save adder
        csa_i: component carry_save_adder
            generic map (
                N => CURRENT_CSA_WIDTH
            )

            port map (
                a  => a_i,
                b  => b_i,
                c  => c_i,
                ps => ps_i,
                cv => cv_i
            );

        -- Extend the partial sum
        ext_ps: component extender
            generic map (
                N_IN            => CURRENT_CSA_WIDTH,
                N_OUT           => CURRENT_CSA_WIDTH + 1,
                TWOS_COMPLEMENT => TWOS_COMPLEMENT
            )

            port map (
                data_in  => ps_i,
                data_out => recursive_signals(WIRE_OFFSETS(IDX_PS + 1) - 1 downto WIRE_OFFSETS(IDX_PS))
            );

        -- Shift the carry vector
        recursive_signals(WIRE_OFFSETS(IDX_CV + 1) - 1 downto WIRE_OFFSETS(IDX_CV)) <= cv_i & '0';
    end generate csa;

    -- TODO: Final ripple carry adder
    sum <= (others => '0');

end architecture behavioral;
